module FourBitAdder(input [3:0] in1, in2, input carry_in, output [3:0] sum, output carry_out);

endmodule